--fil for CTRL