--fil for TX