--fil for CTRL
--test for å se at det fungerer